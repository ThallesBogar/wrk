-- Automatically generated VHDL-93
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use work.all;
use work.mealy_types.all;

entity mealy_topentity_0 is
  port(w3              : in mealy_types.tup2;
       -- clock
       system1000      : in std_logic;
       -- asynchronous reset: active low
       system1000_rstn : in std_logic;
       result          : out signed(8 downto 0));
end;

architecture structural of mealy_topentity_0 is
begin
  mealy_mealy_result : entity mealy_mealy
    port map
      (result          => result
      ,system1000      => system1000
      ,system1000_rstn => system1000_rstn
      ,w2              => w3);
end;
